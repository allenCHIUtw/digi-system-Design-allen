module asu_gate (x, y, mode, carry, out);
input [7:0] x, y;
input mode;
output carry;
output [7:0] out;

/*Write your code here*/
adder_gate the_adder();
barrel_shifter_gate the_shifter();


/*End of code*/


endmodule

module controler(karry,out,md,add,brr);
input
endmodule